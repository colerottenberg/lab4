LIBRARY IeEE; use IeEe.stD_LOgIc_1164.ALl; enTitY FSm IS PoRT ( iD_S_B88665f_7E7082E6_E 
: iN STD_logic; ID_s_b88A71e_7e341cF6_e : In StD_LOgiC; iD_S_5977fb_7FFCC7f4_e : 
in StD_loGic; ID_S_7c95Cc2B_1b9F1D82_E : out stD_logIC; id_S_7c9B02c5_598FA886_e 
: oUT StD_LOgIC; iD_s_34B84a16_43f520dd_E : out stD_lOgIc; iD_S_4BC1c7A7_6B4B6d0F_E 
: oUt stD_LoGIC; id_s_7cA07E8f_1cBd60fa_E : OuT StD_loGIc; ID_S_10B08b40_41C21917_E 
: Out STD_loGIc; iD_S_7cA10aF0_3CF54137_E : OUT STd_LogIC; id_s_10c2A3C1_4193da63_e 
: OUt Std_loGiC; ID_s_7C9844E0_38774De5_e : oUt std_LOgIC; Id_s_fA11bB1_487fE2B_e 
: OUt sTD_loGIC; Id_S_f66e137_35341610_e : iN Std_lOgIc; Id_S_3c0b9Eb_239711A1_E 
: In sTd_logic ); eNd fSm; ARCHItEcTUrE Id_S_5DcFF587_1295F637_E OF FSm Is type iD_S_2DdbF039_4e33D1aa_e 
is (id_S_106149D3_35F88610_e, Id_S_7c988539_38B28d81_E, Id_s_73D8EAE2_7D643Ef5_e, 
iD_S_38d55f9d_45375dC2_E, iD_s_38D55F9e_45375DC3_E, iD_s_19ebFBbB_3A6d6166_E, id_S_19F178e7_266D8Fb4_e, 
iD_S_4012ef9E_5284e514_e, iD_s_3F29fc8a_7f27E122_E); SIgNAl id_S_2DdbF037_4E33d1ac_e, 
id_s_6D8C7f64_12D7C136_E : iD_s_2dDBF039_4E33d1Aa_e; beGin pROcESS(Id_S_B88665f_7e7082E6_e, 
ID_S_B88A71e_7e341Cf6_e) BEgIN If (ID_S_b88a71E_7E341cF6_E = '1') tHeN iD_S_2DdBf037_4e33D1ac_e 
<= id_S_106149d3_35f88610_e; ElsIf (rISInG_EDgE(id_s_b88665f_7e7082E6_e)) Then ID_s_2dDBf037_4e33D1ac_e 
<= ID_S_6d8c7f64_12D7C136_E; EnD if; enD process; PRoCEss(iD_s_5977FB_7ffCC7f4_E, 
ID_S_f66e137_35341610_e, iD_s_3c0B9eb_239711a1_E, iD_s_2DDbf037_4e33D1Ac_e) BeGiN 
id_S_7c95CC2b_1B9f1D82_E <= '0'; iD_s_7c9b02c5_598Fa886_e <= '0'; iD_S_34B84a16_43f520DD_e 
<= '0'; iD_S_4Bc1c7A7_6b4B6d0F_E <= '0'; iD_S_7cA07E8f_1Cbd60Fa_E <= '0'; id_S_10B08B40_41C21917_E 
<= '0'; id_S_7CA10AF0_3cF54137_E <= '0'; Id_s_10c2A3C1_4193dA63_e <= '0'; Id_s_7c9844E0_38774DE5_e 
<= '0'; iD_s_fa11bb1_487fE2b_E <= '0'; iD_S_6D8c7F64_12D7c136_E <= id_s_2ddbf037_4E33D1aC_e;
 CaSe (Id_s_2dDbF037_4e33d1ac_e) IS wHeN id_s_106149d3_35F88610_E => Id_S_7C95cc2b_1B9F1d82_e 
<= '0'; iD_S_4bc1C7A7_6B4B6D0f_e <= '1'; Id_s_34B84A16_43F520dd_e <= '1'; IF (iD_s_5977fB_7ffcC7F4_e 
= '0') ThEN ID_s_6d8C7f64_12d7c136_e <= iD_S_106149d3_35f88610_E; elSE iD_S_6d8c7f64_12d7c136_e 
<= ID_s_7C988539_38b28D81_e; enD If; wHEN Id_S_7C988539_38B28D81_E => iD_s_7C9b02C5_598fA886_E 
<= '1'; iD_s_10B08b40_41C21917_e <= '1'; id_S_7ca07E8f_1cBD60fA_e <= '1'; ID_s_10c2A3c1_4193Da63_e 
<= '1'; ID_S_7ca10aF0_3cf54137_e <= '1'; ID_S_fa11bB1_487Fe2B_E <= '1'; id_S_7C9844E0_38774de5_E 
<= '1'; id_s_7C95cC2b_1B9F1d82_E <= '0'; ID_S_6D8C7f64_12D7c136_E <= ID_S_73d8Eae2_7D643eF5_E;
 when iD_S_73D8eaE2_7d643ef5_e => iF (Id_s_F66e137_35341610_E = '1') thEn ID_S_6D8C7f64_12d7c136_E 
<= iD_S_38D55F9D_45375Dc2_E; ElSE ID_s_6d8C7F64_12d7C136_e <= ID_s_19EBfbbB_3a6D6166_E;
 END If; whEN ID_S_19eBFBbB_3A6D6166_e => If (Id_s_3c0b9eb_239711a1_E = '1') ThEn 
ID_S_6d8c7F64_12D7c136_e <= Id_s_19F178e7_266d8FB4_e; Else Id_s_6D8c7F64_12d7C136_e 
<= ID_S_38D55f9e_45375Dc3_e; EnD if; WHeN id_S_19f178e7_266D8Fb4_e => id_S_10b08B40_41C21917_e 
<= '0'; iD_s_7Ca07e8F_1Cbd60fA_e <= '1'; ID_S_10C2a3c1_4193dA63_E <= '0'; id_S_7CA10AF0_3cF54137_E 
<= '1'; ID_S_fA11bb1_487fe2B_e <= '0'; id_s_7c9844e0_38774DE5_E <= '1'; iD_s_6d8c7f64_12D7C136_E 
<= ID_S_19eBFBBb_3A6d6166_e; wHEn ID_S_38d55f9d_45375dC2_E => id_s_4bC1C7A7_6b4b6d0f_e 
<= '1'; id_S_34B84A16_43f520dD_e <= '1'; id_s_6d8c7f64_12d7c136_E <= id_S_4012Ef9E_5284e514_e;
 wheN Id_S_38D55F9E_45375DC3_e => Id_s_4Bc1C7a7_6b4b6D0f_E <= '0'; Id_s_34B84A16_43f520DD_E 
<= '1'; iD_S_6d8C7F64_12D7c136_e <= ID_s_4012EF9E_5284e514_E; wheN ID_S_4012Ef9E_5284e514_e 
=> iD_s_7c95cc2b_1b9f1d82_e <= '1'; If (iD_s_5977fb_7FFCC7f4_E = '1') theN id_S_6d8c7f64_12D7c136_E 
<= iD_s_4012ef9E_5284e514_e; ELSE iD_S_6D8C7f64_12d7C136_E <= id_s_3F29fc8a_7f27E122_E;
 enD If; when ID_S_3f29Fc8A_7F27e122_e => ID_S_7C95CC2b_1B9F1d82_E <= '1'; If (Id_S_5977Fb_7FFcc7f4_e 
= '0') thEn ID_S_6d8c7f64_12D7c136_E <= ID_S_3F29Fc8a_7F27E122_e; ELSe iD_s_6D8c7F64_12D7C136_e 
<= id_s_7c988539_38b28D81_E; End If; wHeN OtHeRs => null; enD Case; ENd PROCesS; 
eNd id_s_5dcFF587_1295f637_E; 
--------------------------------------------------------------------------------
-- This file was obfuscated and reformated using vHDL Obfuscator GUI          --
-- (c) Miguel Risco-Castillo                                                  --
--------------------------------------------------------------------------------
